module DFlipFlop (clk,A,B);
    input clk, A;
    output B;

    assign B=A;
    
endmodule